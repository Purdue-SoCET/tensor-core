module gsau_top #(
    parameters
) (
    ports
);
    
endmodule