module test_module_tb (
    
);
    test_module test();
endmodule