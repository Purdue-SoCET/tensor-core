module gsau_control_unit #(
    parameters
) (
    ports
);
    
endmodule