`timescale 1ns / 1ns

module benes_tb;
    localparam int PERIOD = 10;
    localparam int SIZE = 32;
    localparam int DWIDTH = 16;
    localparam int TAGWIDTH = $clog2(SIZE);
    localparam int STAGES = (2 * TAGWIDTH) - 1;
    localparam int BITWIDTH = STAGES * (SIZE >> 1);

    logic clk, n_rst;
    logic [BITWIDTH-1:0] control_bit ;

    initial clk = 1'b0;
    always  #5 clk = ~clk;
    
    xbar_if #(.SIZE(SIZE), .DWIDTH(DWIDTH)) xif (.clk(clk), .n_rst(n_rst));
    benes #(.SIZE(SIZE), .DWIDTH(DWIDTH)) DUT (xif, control_bit);

    integer i;
    logic [15:0] val;
    logic [DWIDTH-1:0] exp_out [SIZE-1:0];

    // REQUIRED FOR TESTING WITH CBG

    // typedef logic [DWIDTH-1:0] vec_t [SIZE];
    // vec_t in, exp_out;

    // function automatic void make_vec(output logic [TAGW-1:0] exp_out [SIZE-1:0]);
    //     logic [DWIDTH-1:0] idx [SIZE-1:0];
    //     logic [DWIDTH-1:0] tmp;
    //     integer i, j, tmp;

    //     for (i = 0; i < 32; i++)
    //     idx[i] = i;

    //     for (i = 31; i > 0; i--) begin
    //         j = $urandom_range(0, i); // random index to swap
    //         tmp = idx[i];
    //         idx[i] = idx[j];
    //         idx[j] = tmp;
    //     end

    //     for (i = 0; i < 32; i++)
    //         exp_out[i] = idx[i];

    // endfunction

initial begin
    n_rst = 0;

    #(PERIOD);

    n_rst = 1;
    val = 16'd0;

    for (i = 0; i < 32; i = i + 1) begin
        xif.in[i] = val;
        val = val + 16'd1;
    end
    exp_out = {16'd27, 16'd24, 16'd2, 16'd29, 16'd4, 16'd7, 16'd20, 16'd10, 16'd1, 16'd0, 16'd8, 16'd9, 16'd3, 16'd13, 16'd16, 16'd26,
                    16'd12, 16'd31, 16'd17, 16'd19, 16'd28, 16'd18, 16'd23, 16'd30, 16'd5, 16'd15, 16'd6, 16'd21, 16'd11, 16'd25, 16'd22, 16'd14};
    
    control_bit = 144'b111000110101110001100100110011100111001110000000111100000001101100101011001100000000000000000000001000011001000001110110011110001011111001001100;  
    
    repeat (10) #(PERIOD);
    
    for (i = 0; i < 32; i = i + 1) begin
        if(xif.out[i] != exp_out[(SIZE-1 - i)]) begin
            $display("wrong output for %d", i);
        end
        // $display("output %d: %d", i, xif.out[i]);
    end
    $finish;
end

endmodule












`timescale 1ns/1ns

`include "xbar_params.svh"
`include "xbar_if.sv"
`include "cbg_benes.sv"

module benes_tb;

  import xbar_pkg::*;

  localparam int SIZE = 32;
  localparam int DWIDTH = 16;
  localparam int TAGW = $clog2(SIZE);
  localparam int STAGES = (2 * TAGW) - 1; // 9 for SIZE=32
  localparam int BITWIDTH = STAGES * (SIZE >> 1); // 9 * 16 = 144
  localparam logic [STAGES-2:0] REGISTER_MASK = 8'b11111111;
  localparam int REAL_LATENCY = $countones(REGISTER_MASK) + 1;
  localparam int N_REQS = (REAL_LATENCY * 2);
  localparam int VERBOSE = 0;
  localparam bit PERM_IS_OUT_TO_IN = 1;

  logic clk, n_rst;
  initial clk = 1'b0;
  always #5 clk = ~clk;

  xbar_if #(.SIZE(SIZE), .DWIDTH(DWIDTH)) xif (.clk(clk), .n_rst(n_rst));

  logic [BITWIDTH-1:0] control_bit;

  benes #(.SIZE(SIZE), .DWIDTH(DWIDTH), .REGISTER_MASK(REGISTER_MASK)) dut (.xif(xif.xbar), .control_bit(control_bit));

  logic [TAGW-1:0] perm_cfg [SIZE]; // feed to CBG
  logic [BITWIDTH-1:0] ctrl; // control bits produced by CBG

  cbg_benes #(.SIZE(SIZE)) cbg (.perm(perm_cfg), .ctrl(ctrl));

  typedef logic [DWIDTH-1:0] vec_t [SIZE];
  vec_t exp_q[$]; // queue of expected vectors 

  // Fill with randome values
  function automatic void make_vec(output vec_t v);
    for (int i = 0; i < SIZE; i++) v[i] = $urandom();
  endfunction

  // OUT->IN permutation generator using Fisher–Yates:
  // out_to_in[o] = index of input that should appear at output o
  function automatic void make_random_perm_out_to_in(output logic [TAGW-1:0] out_to_in [SIZE]);
    int idx [SIZE];
    for (int i = 0; i < SIZE; i++) begin 
        idx[i] = i;
    end
    for (int k = SIZE-1; k > 0; k--) begin
      int j = $urandom_range(0, k);
      int t = idx[k]; idx[k] = idx[j]; idx[j] = t;
    end
    for (int o = 0; o < SIZE; o++) begin 
        out_to_in[o] = TAGW'(idx[o]);
    end
  endfunction

  // If p_out_in[o] = i, produce p_in_out[i] = o
  function automatic void invert_perm(input  logic [TAGW-1:0] p_out_in [SIZE], output logic [TAGW-1:0] p_in_out [SIZE]);
    for (int i = 0; i < SIZE; i++) begin 
        p_in_out[i] = 'x;
    end
    for (int o = 0; o < SIZE; o++) begin 
        p_in_out[p_out_in[o]] = TAGW'(o);
    end
  endfunction

  // Apply OUT->IN permutation to form expected: exp[o] = in[p[o]]
  function automatic void apply_perm_o2i(input vec_t in_vec, input logic [TAGW-1:0] p [SIZE], output vec_t exp);
    for (int o = 0; o < SIZE; o++) begin 
        exp[o] = in_vec[p[o]];
    end
  endfunction

  int launched, retired, errors;
  int mismatches;

  initial begin : main
    vec_t in_vec, exp_vec, exp;
    logic [TAGW-1:0] perm_out_to_in [SIZE];
    logic [TAGW-1:0] perm_in_to_out [SIZE];
    logic [DWIDTH-1:0] got;

    n_rst = 1'b0;
    xif.en = 1'b0;
    control_bit = '0;
    for (int i = 0; i < SIZE; i++) begin
      xif.in[i].din   = '0;
      xif.in[i].shift = TAGW'(i); 
    end
    repeat (5) @(posedge clk);
    n_rst = 1'b1;
    @(posedge clk);

    // 1 permutation for the whole streaming window (control held steady)
    make_random_perm_out_to_in(perm_out_to_in);

    // permutation into CBG 
    if (PERM_IS_OUT_TO_IN) begin
      for (int i = 0; i < SIZE; i++) begin 
        perm_cfg[i] = perm_out_to_in[i];
      end
    end else begin
      invert_perm(perm_out_to_in, perm_in_to_out);
      for (int i = 0; i < SIZE; i++) begin
        perm_cfg[i] = perm_in_to_out[i];
      end
    end

    control_bit = ctrl;
    launched = 0;
    retired  = 0;
    errors   = 0;
    xif.en = 1'b1;

    for (int t = 0; t < N_REQS; t++) begin
      if (launched <= REAL_LATENCY) begin
        make_vec(in_vec);
        apply_perm_o2i(in_vec, perm_out_to_in, exp_vec);
        exp_q.push_back(exp_vec);
        launched++;
        // Drive one full vector 
        for (int i = 0; i < SIZE; i++) begin
          xif.in[i].din   = in_vec[i];
          xif.in[i].shift = TAGW'(i);
        end
      end

      @(posedge clk);
      if (launched >= REAL_LATENCY) begin
        exp = exp_q.pop_front();
        mismatches = 0;

        for (int k = 0; k < SIZE; k++) begin
          got = xif.out[k];
          if (got !== exp[k]) begin
            mismatches++;
            errors++;
            $display($sformatf("[BENES][lane%0d] got=%0d exp=%0d", k, got, exp[k]));
          end else if (VERBOSE) begin
            $display($sformatf("[BENES][lane%0d] got=%0d exp=%0d", k, got, exp[k]));
          end
        end

        if (mismatches == 0) begin
          $display("[BENES][Complete] retire=%0d OK", retired);
        end else begin
          $display("[BENES][Complete] retire=%0d mismatches=%0d", retired, mismatches);
        end
        retired++;
      end
    end

    xif.en = 1'b0;
    $display("[BENES][Summary] errors=%0d (latency=%0d)", errors, REAL_LATENCY);
    $finish;
  end

endmodule
