`include "scpad_types_pkg.vh"
`include "scratchpad_if.vh"

module frontend (
    input logic clk, n_rst,
    scpad_if.frontend fcif
); 
    import scpad_types_pkg::*;


endmodule