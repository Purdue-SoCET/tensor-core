`ifndef SOCETLIB_COUNTER_IF
`define SOCETLIB_COUNTER_IF


`endif