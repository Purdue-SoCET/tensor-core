module test_module(
    
);
    
endmodule