module sqrt_pipe_tb;


endmodule