module param_sr_tb;


endmodule