/*  Haejune Kwon - kwon196@purdue.edu */
/*  Akshath Raghav Ravikiran - araviki@purdue.edu */

`include "xbar_params.svh"
`include "xbar_if.sv"

module benes_xbar #(
    parameter int SIZE = 32,
    parameter int DWIDTH = 16
) (xbar_if.xbar xif);

endmodule