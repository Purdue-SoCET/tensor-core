`include "scpad_types_pkg.vh"
`include "scratchpad_if.vh"

module xbar (
    input logic clk, n_rst,
    scpad_if.xbar xif
); 
    import scpad_types_pkg::*;

endmodule