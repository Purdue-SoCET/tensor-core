`ifndef  SCRATCHPAD_IF_VH
`define SCRATCHPAD_IF_VH
`include "types_pkg.vh"

interface scratchpad_if;
    import types_pkg::*;
    
    

    modport sp (
        input 
        output 
    );
    

endinterface

`endif 