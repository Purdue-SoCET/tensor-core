`ifndef XBAR_PARAMS_SVH
`define XBAR_PARAMS_SVH

    parameter int unsigned NAIVE_LATENCY   = 1;
    parameter int unsigned BENES_LATENCY   = 3;
    parameter int unsigned BATCHER_LATENCY = 4;
    
`endif
