`ifndef DRAM_REQ_QUEUE_IF
`define DRAM_REQ_QUEUE_IF

`include "scpad_pkg.sv"
`include "scpad_if.sv"

interface dram_req_queue_if;
    import scpad_pkg::*;

    logic sched_write;
    dram_req_t dram_req;
    logic [DRAM_ADDR_WIDTH-1:0] dram_addr;
    logic [DRAM_ID_WIDTH-1:0]   id;
    logic [2:0]   sub_id, num_request;
    logic [DRAM_VECTOR_MASK-1:0]   dram_vector_mask;
    scpad_data_t sram_rdata;
    logic be_stall, sched_valid;
    logic dram_queue_full, dram_be_stall, sram_res_valid, burst_complete;
    logic transaction_complete, initial_request_done;

    modport baceknd_dram_req_queue ( 
        input dram_addr, id, sub_id, dram_vector_mask, sram_rdata, sram_res_valid, num_request, sched_valid,
        input sched_write,       // scheduler write = 1 means it's a scpad store aka we need to do a dram write.
        input be_stall, initial_request_done,
        input dram_be_stall,     // tells us if the dram is ready to accept our req. If it is and our FIFO is valid then we can assume 
                                  // our current req will be successfully latched in the dram controller and can invalidate nxt cycle
        output dram_req, dram_queue_full, burst_complete, transaction_complete
    );

endinterface

`endif //DRAM_REQ_QUEUE_IF