module gsau_queue #(
    parameters
) (
    ports
);
    
endmodule