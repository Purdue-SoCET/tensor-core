`include "scpad_types_pkg.vh"
`include "scratchpad_if.vh"

module backend (
    input logic clk, n_rst,
    scpad_if.backend bif
); 

endmodule