`include "scratchpad_if.vh"

module scratchpad ()