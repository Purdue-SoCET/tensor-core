import scpad_pkg::*;

module backend #(parameter logic [SCPAD_ID_WIDTH-1:0] IDX = '0) (scpad_if.backend_sched bshif, scpad_if.backend_scpads bscif, scpad_if.backend_dram bdrif); 

    // grab clk and n_rst from any 

endmodule