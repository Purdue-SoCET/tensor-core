`include "scpad_types_pkg.vh"
`include "scratchpad_if.vh"

module frontend_vc (
    input logic clk, n_rst,
    scpad_if.frontend fif
); 
    import scpad_types_pkg::*;

endmodule