`include "swizzle_if.vh"
import scpad_pkg::*;

module swizzle (
  swizzle_if.swizzle sw
);

    logic [ROW_IDX_WIDTH-1:0] abs_row;

    always_comb begin
        sw.xbar_desc.valid_mask = '0;
        sw.xbar_desc.shift_mask = '0;
        sw.xbar_desc.slot_mask  = '0;

        for (int bank_id = 0; bank_id < NUM_COLS; bank_id++) begin
            if (sw.row_or_col) begin // row-major read
                abs_row = sw.spad_addr + sw.row_id;
                sw.xbar_desc.valid_mask[bank_id] = (bank_id < sw.num_cols);
                sw.xbar_desc.shift_mask[bank_id] = COL_IDX_WIDTH'((bank_id ^ (abs_row & (NUM_COLS-1))) & (NUM_COLS-1));
                sw.xbar_desc.slot_mask[bank_id]  = abs_row;
            end else begin
                abs_row = base_row + ROW_IDX_WIDTH'(bank_id);
                sw.xbar_desc.valid_mask[bank_id] = (bank_id < sw.num_rows);
                sw.xbar_desc.shift_mask[bank_id] = COL_IDX_WIDTH'((sw.col_id ^ (abs_row & (NUM_COLS-1))) & (NUM_COLS-1));
                sw.xbar_desc.slot_mask[bank_id]  = abs_row;
            end
        end
    end

endmodule


