`ifndef DRAM_TOP_VH
`define DRAM_TOP_VH
`include "dram_pkg.vh"


interface dram_top_if();


    

endinterface

`endif